//READ ONLY VEDA MEMORY
module instrMemory (
	input clk,
	input  [ 5:0] addr,
	output [31:0] data
);

	reg [31:0] data;
	reg [31:0] memory [63:0];

	initial begin
		
			//jumps to bubbel sort execution, skipping the test instructions
			memory[0] = 32'b000111_000000_000000_000000_00001001; //j #04
		
			//test instructions: to check each instruction used in bubble sort
			memory[1] = 32'b000001_00000_00010_0000000000000101; //addi $2, $0, 5
			memory[2] = 32'b000001_00000_00011_0000000000000101; //addi $3, $0, 3
			memory[3] = 32'b000000_00010_00011_00100_00000_000000; //add $4, $2, $3
			memory[4] = 32'b000010_00100_00101_0000000000000010; //sll $5, $4, 2
			memory[5] = 32'b000011_00100_00101_00110_00000_000000; //slt $6, $5, $4
			memory[6] = 32'b000100_00000_00101_0000000000000000; //sw $5, (0)$zero
			memory[7] = 32'b000101_00000_00110_0000000000000000; //lw $6, (0)$zero
			memory[8] = 32'b000110_00010_00011_0000000000000001; //beq $2, $3, #04

			//bubble sort machine code
			memory[9] = 32'b000001_00000_00001_0000000000000000; //li $s0, 0
			memory[10] = 32'b000101_00000_00111_0000000000000001; //lw $s6, N-1;
			memory[11] = 32'b000101_00000_01110_0000000000000000; //lw $t4, N;
			memory[12]= 32'b000001_00000_01101_0000000000000000; //li $t3, 0;
			memory[13] = 32'b000001_00000_00010_0000000000000000; //li $s1, 0;
			memory[14] = 32'b000001_00000_01000_0000000000000010; //la $s7, numbers;
			memory[15] = 32'b000001_00010_10001_0000000000000000; //sll $t7, $s1, 0;
			memory[16] = 32'b000000_10001_01000_10001_00000_000000; //add $t7, $s7, $t7 
			memory[17] = 32'b000101_10001_01010_0000000000000000; //lw $t0, 0($t7)  
			memory[18] = 32'b000101_10001_01011_0000000000000001; //lw $t1, 4($t7)
			memory[19] = 32'b000011_01010_01011_01100_00000_000000; //slt $t2, $t0, $t1	
			memory[20] = 32'b000110_00000_01100_0000000000000001; //beq $t2, $zero, swap
			memory[21] = 32'b000111_000000_000000_000000_00011000; //j increment
			memory[22] = 32'b000100_10001_01011_0000000000000000; //sw $t1, 0($t7) 
			memory[23] = 32'b000100_10001_01010_0000000000000001; //sw $t0, 4($t7)
			memory[24] = 32'b000001_00010_00010_0000000000000001; //	addi $s1, $s1, 1				
			memory[25] = 32'b000000_00010_00001_00110_00000_000000; //add $s5, $s1, $s0 	
			memory[26] = 32'b000110_00111_00110_0000000000000001; //beq $s6, $s5, continue
			memory[27] = 32'b000111_000000_000000_000000_00001111; //j loop
			memory[28] = 32'b000001_00001_00001_0000000000000001; //addi $s0, $s0, 1
			memory[29] = 32'b000001_00000_00010_0000000000000000; //li $s1, 0
			memory[30] = 32'b000110_00001_00111_0000000000000001; //beq $s0, $s6, continue
			memory[31] = 32'b000111_000000_000000_000000_00001111; //j loop

			// memory[32] = 32'b000101_00000_01010_0000000000000000;
			// memory[33] = 32'b000101_00000_01010_0000000000000001;
			
			//data memory is now filled with the sorted array
			memory[32] = 32'b000101_00000_01010_0000000000000010;
			memory[33] = 32'b000101_00000_01010_0000000000000011;
			memory[34] = 32'b000101_00000_01010_0000000000000100;
			memory[35] = 32'b000101_00000_01010_0000000000000101;
			memory[36] = 32'b000101_00000_01010_0000000000000110;
			memory[37] = 32'b000101_00000_01010_0000000000000111;
			memory[38] = 32'b000101_00000_01010_0000000000001000;
			memory[39] = 32'b000101_00000_01010_0000000000001001;
			memory[40] = 32'b000101_00000_01010_0000000000001010;

			memory[41] = 32'h00000000;
			memory[42] = 32'h00000000;
			memory[43] = 32'h00000000;
			memory[44] = 32'h00000000;
			memory[45] = 32'h00000000;
			memory[46] = 32'h00000000;
			memory[47] = 32'h00000000;
			memory[48] = 32'h00000000;
			memory[49] = 32'h00000000;
			memory[50] = 32'h00000000;
			memory[51] = 32'h00000000;
			memory[52] = 32'h00000000;
			memory[53] = 32'h00000000;
			memory[54] = 32'h00000000;
			memory[55] = 32'h00000000;
			memory[56] = 32'h00000000;
			memory[57] = 32'h00000000;
			memory[58] = 32'h00000000;
			memory[59] = 32'h00000000;
			memory[60] = 32'h00000000;
			memory[61] = 32'h00000000;
			memory[62] = 32'h00000000;
			memory[63] = 32'h00000000;
	end

	always @(*) begin
		data = memory[addr];
	end

endmodule
